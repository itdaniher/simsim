* AD8018 Spice Model
* Description: Amplifier
* Generic Desc: Dual 350mA 135MHz high output drivers
* Developed by: BJG
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (09/2000)
* Copyright 2000, 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement.
* Use of this model indicates your acceptance with the terms and provisions in the License Statement
*
* BEGIN Notes:
*
* Not Modeled:
*       Eref is not refered to ground, rather it is set to a point midway between supply voltages
*       distortion is not characterized
*
* Parameters modeled include:
*       open loop gain and phase vs. frequency (modeled to fit performance with 5 ohm load and to maintain stability
*       output clamping voltage and current
*	Input offset voltage and bias currents
*       slew rate
*       output currents are reflected to V supplies
*
* END Notes
*
* Node assignments
*                   non-inverting input
*                   | inverting input
*                   | | positive supply
*                   | | |  negative supply
*                   | | |  |  output
*                   | | |  |  |
.subckt AD8018      3 2 7  4  1

***** Input stage ********
Q1         7 31 210 QN
Q2         4 31 156 QP
Q3         670 156 196 QN
Q4         665 210 196 QP
I1         210 4 DC 1.04e-4
I2         7 156 DC 1.04e-4
R1         7 670  1k
R2         665 4  1k
C2         3 4  .5e-18
C5         2 7  .35e-12
C6         4 2  .35e-12
L2         196 2 1nH

***** Input Error Sources *****
EOS         31 3 POLY(1) 643 100 (1.804e-3,1)
GB1         7 3 POLY(1) 3 100 (1e-6,1e-15)
GB2         7 2 POLY(1) 3 100 (0.6e-6,1e-15)


***** Reference Stage
EREF         100 0 POLY(2) (7,0) (4,0) (0,.5,.5)


***** Gain Stage *****
D1         6048 670 diode
D2         665 6102 diode
V1         7 6048 DC .47
V2         6102 4 DC .47
G1         100 1569 7 670 0.118e-3
G2         1569 100 665 4 0.118e-3
R3         1569 100 21000k
C1         1569 100 .37e-12

D3         1569 1721 diode
D4         1747 1569 diode
VOC1       7 1721 1.08
VOC2       1747 4 1.05


***** CMRR Stage *****

ECM         100 1977 3 100 19.95
CCM         1977 643  3.68e-11
RCM1         1977 643  500
RCM2         643 100  1


***** Pole at 100 MHz  *****

G4         100 319 6844 100 1e-6
C4         100 319 1.59e-15
R5         100 319 1000k


***** Pole at 600 MHz +*****

G3         100 6844 1569 100 1e-6
R4         100 6844  1000k
C3         100 6844  .265e-15


*****Output Stage *****

VW         319 268 DC 0

DSC1         268 2713 diode
DSC2         2716 268 diode
VSC1         2713 2751 DC -.3
VSC2         2751 2716 DC -.3

DSY1         313 314 diode
DSY2         315 313 diode
VSY1         314 100 DC 0
VSY2         100 315 DC 0
GSY         100 313 2751 268 10

GO1         2751 7 7 268 10
GO2         4 2751 268 4 10
RO1         7 2751  .1
RO2         2751 4  .1
L1         2751 1  1nH
FSY         7 4 POLY(2) VSY1 VSY2 8.699E-3 1 1


.model diode D (IS=10E-15)
.model QN NPN (Is=2.57e-17 Bf=110 Vaf=100)
.model QP PNP (Is=2.49e-17 Bf=93 Vaf=23.8)
.ends





