* ADA4661-2 SPICE Macro-model
* Typical Values
* 07/13, Version 0
* VW ADSJ
*
* Copyright 2013 by Analog Devices
*
* VSY=18V, T=25�C
*
* Refer to "README.DOC" file for License Statement.  Use of this
* model indicates your acceptance of the terms and provisions in
* the License Statement.
*
* Node Assignments
*                       noninverting input
*                       |   inverting input
*                       |   |    positive supply
*                       |   |    |   negative supply
*                       |   |    |   |   output
*                       |   |    |   |   |
*                       |   |    |   |   |
.SUBCKT ADA4661         1   2   99  50  45
*
* INPUT STAGE
*
M1   4  7  8  8 PIX L=1E-6 W=2.65E-04
M2   6  2  8  8 PIX L=1E-6 W=2.65E-04
M3  14  7 18 18 NIX L=1E-6 W=1.18E-04
M4  16  2 18 18 NIX L=1E-6 W=1.18E-04
RD1  4 50 1.33E+04
RD2  6 50 1.33E+04
RD3 99 14 1.33E+04
RD4 99 16 1.33E+04
C1   4  6 8.15E-13
C2  14 16 8.15E-13
I1  99  8 3.00E-05
I2  18 50 3.00E-05
V1  99  9 2.113E+00 
V2  19 50 1.203E-01 
D1   8  9 DX
D2  19 18 DX
EOS  7  1 POLY(4) (73,98) (22,98) (81,98) (83,98) 1.50E-04 1 1 1 1
IOS  1  2 1.50E-12
Ccm1 1 50 3E-12
Ccm2 2 50 3E-12
Cdm 1 2 8.5E-12
*
*CMRR
*
E1  72 98 POLY(2) (1,98) (2,98) 0 5.25E-03 5.25E-03
R10 72 73 1.89E+02
R20 73 98 7.959E-02
C10 72 73 1.00E-06
*
* PSRR
*
EPSY 21 98 POLY(1) (99,50) -2.074E+02 1.152E+1
RPS1 21 22 1.59E+05
RPS2 22 98 3.18E-02
CPS1 21 22 1.00E-06
*
* VOLTAGE NOISE 
*
VN1 80 98 0
RN1 80 98 16.45E-3
HN  81 98 VN1 1.07E+01
RN2 81 98 1
*
* FLICKER NOISE CORNER 
*
DFN 82 98 DNOISE
VFN 82 98 DC 0.6441
HFN 83 98 POLY(1) VFN 1.00E-03 1.00E+00
RFN 83 98 1
*
* INTERNAL VOLTAGE REFERENCE
*
EREF 98  0 POLY(2) (99,0) (50,0) 0 0.5 0.5
GSY  99 50 POLY(1) (99,50) 4.575E-04 -1.55E-6
EVP  97 98 POLY(1)(99,50) 0.5 0.175
EVN  51 98 POLY(1)(50,99) 0.5 0.375
*
* GAIN STAGE
*
G1 98 30 POLY(2) (4,6) (14,16) 0 7.103E-03 7.103E-03
R1 30 98 1.00E+06
RZ 455 31 0.195E+00
CF 30 31 2.95E-9
EZ 455 98 (45,98) 1
D3 30 97 DX
D4 51 30 DX
*
* OUTPUT STAGE
*
M5  45 46 99 99 POX L=3E-6 W=5.99E-04
M6  45 47 50 50 NOX L=3E-6 W=5.99E-03
EG1 99 46 POLY(1) (98,30) 8.523E-01 1
EG2 47 50 POLY(1) (30,98) 6.964E-01 1

*
* MODELS
*
.MODEL POX PMOS (LEVEL=2,KP=4.00E-05,VTO=-0.7,LAMBDA=0.047,RD=0)
.MODEL NOX NMOS (LEVEL=2,KP=1.00E-05,VTO=+0.6,LAMBDA=0.022,RD=0)
.MODEL PIX PMOS (LEVEL=2,KP=1.50E-05,VTO=-0.5,LAMBDA=0.047)
.MODEL NIX NMOS (LEVEL=2,KP=4.00E-05,VTO=0.5,LAMBDA=0.022)
.MODEL DX D(IS=1E-14,RS=0.1)
.MODEL DNOISE D(IS=1E-14,RS=0,KF=1.53E-10)
*
*
.ENDS ADA4661
*
*$
