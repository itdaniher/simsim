.TITLE "ada4661 test"

.INCLUDE ./models/ada4661.cir

X4661 ni ii vss vdd vo ADA4661

VS vdd vss DC 7
VGND vdd vgnd DC 1

VIN vgnd ni DC 2.5 AC 1

Rf ii vo 0
Rl vo vgnd 100

.control
tf v(vo,ni) vin
print all
ac dec 10 10 100meg
plot v(vo)
plot phase(v(vo))
.endc
.end
